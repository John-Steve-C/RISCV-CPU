module RS(

);

endmodule