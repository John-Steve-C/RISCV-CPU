module ALU(
    input wire clk_in,
    input wire rst_in
);



endmodule