module RoB(

);

endmodule