module ALU(
    input wire clk_in,
    input wire rst_in,

    input wire [31:0] rs1,
    input wire [31:0] rs2,
    input wire [31:0] rd
);



endmodule